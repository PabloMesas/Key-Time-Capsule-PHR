LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

CONSTANT a : INTEGER := 2;

ENTITY MODEXP IS
PORT (t : IN STD_LOGIC_VECTOR(1023 DOWNTO 0);
      n : IN STD_LOGIC_VECTOR(1024 DOWNTO 0);
      s : OUT STD_LOGIC_VECTOR(1023 DOWNTO 0);
     );
END MODEXP;

ARCHITECTURE ARC OF MODEXP IS
  VARIABLE a : IN STD_LOGIC_VECTOR(1024 DOWNTO 0);
  BEGIN
    IF t <= 0 THEN a = 1;
    ELSE
      FOR i in 0 to t loop:
        a sll 1;
	IF a > n THEN
	  a = a - n;
	END IF;
      END LOOP;
    END IF;
END ARC;
