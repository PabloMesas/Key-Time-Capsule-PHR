LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TestPowMod IS
END TestPowMod;

ARCHITECTURE testbasics OF TestPowMod IS

COMPONENT PowerModulus
PORT (a, t, n : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
      r : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
     );
END COMPONENT;

SIGNAL a, t, n, r: STD_LOGIC_VECTOR(127 DOWNTO 0);

BEGIN

I1: PowerModulus PORT MAP (a, t, n, r);

a <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010" after 0 ns,
     "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011" after 20 ns, 
     "00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010" after 40 ns;

t <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101" after 0 ns,
     "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101" after 20 ns, 
     "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011" after 40 ns;

n <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111" after 0 ns,
     "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111" after 20 ns, 
     "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000" after 40 ns;

END testbasics; 